module core (
    
);

endmodule